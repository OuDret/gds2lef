MACRO NAND
	CLASS CORE ;
	ORIGIN 0 0 ;
	FOREIGN NAND 0 0 ;
	SIZE 6.29 BY 5.46 ;
	SYMMETRY X Y ;
	SITE std_cell ;
	OBS 
		LAYER metal2 ;
			RECT -2.46 -1.23 -1.33 3.95 ;
			POLYGON 3.23 -2.45 -0.77 -1.98 -1.09 0.4 1.92 -0.87 1.61 0.56 3.41 2.37 ;
	END
	PIN A
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal3 ;
			RECT -1.77 1.11 -0.51 2.27 ;
	END A
	PIN B
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal3 ;
			RECT 0.6 3.1 1.69 4.33 ;
	END B
	PIN Y
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal3 ;
			RECT 3.87 1.31 5.36 2.8 ;
	END Y
	OBS 
		LAYER via ;
			POLYGON 5.76 -2.67 1.83 2.17 -1.34 3.24 2.14 5.46 5.57 3.66 ;
			POLYGON -1.14 -2.37 -3.09 -1.6 -2.25 -0.53 -0.57 -0.72 ;
	END
END

MACRO NOR
	CLASS CORE ;
	ORIGIN 0 0 ;
	FOREIGN NOR 0 0 ;
	SIZE 25.31 BY 21.95 ;
	SYMMETRY X Y ;
	SITE std_cell ;
	OBS 
		LAYER metal2 ;
			POLYGON 4.99 6.13 0.0 14.08 7.42 21.36 9.98 21.95 9.85 10.14 ;
	END
	OBS 
		LAYER metal3 ;
			POLYGON 10.8 0.0 10.8 1.5 21.55 1.56 21.39 8.04 16.35 7.85 16.34 7.87 16.24 12.84 16.26 12.87 25.31 12.71 25.29 11.21 17.77 11.35 17.8 9.41 22.84 9.6 22.85 9.59 23.09 0.08 23.07 0.06 ;
	END
	PIN A
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER via ;
			RECT 8.51 8.82 11.61 12.05 ;
	END A
	PIN Y
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER via ;
			RECT 15.98 14.91 19.05 19.24 ;
	END Y
	OBS 
		LAYER via ;
			RECT 16.15 2.18 19.98 5.96 ;
	END
END

