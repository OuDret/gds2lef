MACRO NOR
	CLASS CORE ;
	ORIGIN 0 0 ;
	FOREIGN NOR 0 0 ;
	SIZE 131.5 BY 340 ;
	SYMMETRY X Y ;
	SITE std_cell ;
	OBS 
		LAYER metal2 ;
			POLYGON -9.65 1.64 -14.64 9.59 -7.22 16.87 -4.66 17.46 -4.79 5.65 ;
	END
	OBS 
		LAYER metal3 ;
			POLYGON -3.84 -4.49 -3.84 -2.99 6.91 -2.93 6.75 3.55 1.71 3.36 1.7 3.38 1.6 8.35 1.62 8.38 10.67 8.22 10.65 6.72 3.13 6.86 3.16 4.92 8.2 5.11 8.21 5.1 8.45 -4.41 8.43 -4.43 ;
	END
	PIN A
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER via ;
			RECT -6.13 4.33 -3.03 7.56 ;
	END A
	PIN Y
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER via ;
			RECT 1.34 10.42 4.41 14.75 ;
	END Y
	OBS 
		LAYER via ;
			RECT 1.51 -2.31 5.34 1.47 ;
	END
END

MACRO NAND
	CLASS CORE ;
	ORIGIN 0 0 ;
	FOREIGN NAND 0 0 ;
	SIZE 131.5 BY 340 ;
	SYMMETRY X Y ;
	SITE std_cell ;
	OBS 
		LAYER metal2 ;
			RECT -2.46 -1.23 -1.33 3.95 ;
			POLYGON 3.23 -2.45 -0.77 -1.98 -1.09 0.4 1.92 -0.87 1.61 0.56 3.41 2.37 ;
	END
	PIN A
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal3 ;
			RECT -1.77 1.11 -0.51 2.27 ;
	END A
	PIN B
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal3 ;
			RECT 0.6 3.1 1.69 4.33 ;
	END B
	PIN Y
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal3 ;
			RECT 3.87 1.31 5.36 2.8 ;
	END Y
	OBS 
		LAYER via ;
			POLYGON 5.76 -2.67 1.83 2.17 -1.34 3.24 2.14 5.46 5.57 3.66 ;
			POLYGON -1.14 -2.37 -3.09 -1.6 -2.25 -0.53 -0.57 -0.72 ;
	END
END

